magic
tech sky130A
magscale 1 2
timestamp 1739896874
<< error_p >>
rect 4286 8538 4318 8540
rect 4192 7278 4196 7280
rect 4192 7244 4196 7246
rect 5737 4973 5739 4988
rect 5737 4945 5738 4960
rect 27416 492 27420 494
<< error_s >>
rect 15820 41896 15822 41898
rect 15818 41894 15822 41896
rect 15272 41892 15278 41894
rect 15816 41892 15822 41894
rect 15278 41886 15284 41892
rect 15810 41886 15816 41892
rect 5035 41678 5047 41690
rect 5369 41678 5381 41690
rect 5035 41672 5381 41678
rect 5035 41332 5381 41338
rect 5035 41320 5047 41332
rect 5369 41320 5381 41332
rect 5524 5198 5526 5210
rect 5552 5184 5554 5194
<< locali >>
rect 3616 4330 4334 4364
rect 3616 3998 3640 4330
rect 4310 3998 4334 4330
rect 3616 3984 4334 3998
<< viali >>
rect 5035 41332 5381 41678
rect 3640 3998 4310 4330
<< metal1 >>
rect 5025 41332 5035 41678
rect 5381 41332 5391 41678
rect 3606 4002 3616 4354
rect 4324 4002 4334 4354
rect 3616 3998 3640 4002
rect 4310 3998 4330 4002
rect 3616 3984 4330 3998
<< via1 >>
rect 5035 41332 5381 41678
rect 3616 4330 4324 4354
rect 3616 4002 3640 4330
rect 3640 4002 4310 4330
rect 4310 4002 4324 4330
<< metal2 >>
rect 15276 43600 15822 43610
rect 15268 43100 15276 43588
rect 15822 43100 15834 43588
rect 15268 42858 15834 43100
rect 15272 42548 15820 42858
rect 15280 41896 15820 42548
rect 5035 41678 5381 41688
rect 5035 41322 5381 41332
rect 3616 4354 4324 4364
rect 3616 3992 4324 4002
<< via2 >>
rect 15276 43100 15822 43600
rect 5035 41332 5381 41678
rect 3616 4002 4324 4354
<< metal3 >>
rect 15284 43608 15830 43612
rect 15284 43605 27416 43608
rect 15266 43600 27416 43605
rect 15266 43100 15276 43600
rect 15822 43108 27416 43600
rect 15822 43100 15832 43108
rect 15266 43095 15832 43100
rect 5025 41678 5391 41683
rect 782 41328 792 41678
rect 1200 41332 5035 41678
rect 5381 41332 5391 41678
rect 1200 41328 1440 41332
rect 5025 41327 5391 41332
rect 3606 4354 4334 4359
rect 3606 4348 3616 4354
rect 1398 4342 3616 4348
rect 1380 3992 1390 4342
rect 1798 4002 3616 4342
rect 4324 4002 4334 4354
rect 1798 3997 4334 4002
rect 1798 3996 4008 3997
rect 1798 3992 1808 3996
rect 27018 520 27416 43108
rect 27224 492 27416 520
rect 27224 438 27420 492
rect 27224 304 27238 438
rect 27408 434 27420 438
rect 27408 304 27416 434
rect 27224 296 27416 304
<< via3 >>
rect 792 41328 1200 41678
rect 5035 41332 5381 41678
rect 1390 3992 1798 4342
rect 27238 304 27408 438
<< metal4 >>
rect 3006 44952 3066 45152
rect 3558 44952 3618 45152
rect 4110 44952 4170 45152
rect 4662 44952 4722 45152
rect 5214 44952 5274 45152
rect 5766 44952 5826 45152
rect 6318 44952 6378 45152
rect 6870 44952 6930 45152
rect 7422 44952 7482 45152
rect 7974 44952 8034 45152
rect 8526 44952 8586 45152
rect 9078 44952 9138 45152
rect 9630 44952 9690 45152
rect 10182 44952 10242 45152
rect 10734 44952 10794 45152
rect 11286 44952 11346 45152
rect 11838 44952 11898 45152
rect 12390 44952 12450 45152
rect 12942 44952 13002 45152
rect 13494 44952 13554 45152
rect 14046 44952 14106 45152
rect 14598 44952 14658 45152
rect 15150 44952 15210 45152
rect 15702 44952 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 44952 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 200 1000 600 44152
rect 800 41679 1200 44152
rect 791 41678 1201 41679
rect 791 41328 792 41678
rect 1200 41328 1201 41678
rect 791 41327 1201 41328
rect 800 1000 1200 41327
rect 1400 4343 1800 44152
rect 5034 41678 5382 41679
rect 5034 41332 5035 41678
rect 5381 41332 5382 41678
rect 5034 41331 5382 41332
rect 1389 4342 1800 4343
rect 1389 3992 1390 4342
rect 1798 3992 1800 4342
rect 1389 3991 1800 3992
rect 1400 1000 1800 3991
rect 27232 438 27416 450
rect 27232 304 27238 438
rect 27408 304 27416 438
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27232 172 27416 304
rect 27234 0 27414 172
use bandgap  bandgap_0
timestamp 1739894026
transform 0 -1 6280 1 0 634
box 3348 -10162 41804 2662
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
