magic
tech sky130A
magscale 1 2
timestamp 1739894026
<< error_s >>
rect 6610 2084 6612 2088
rect 6644 2084 6646 2088
rect 7904 1962 7906 1994
rect 4564 754 4588 756
rect 4550 726 4560 728
rect 4311 542 4326 543
rect 4339 541 4354 543
rect 41258 -8998 41260 -8992
rect 41252 -9004 41258 -8998
rect 41252 -9536 41258 -9530
rect 41652 -9536 41656 -9530
rect 41258 -9538 41260 -9536
rect 41258 -9542 41264 -9538
rect 41644 -9542 41650 -9538
<< nwell >>
rect 6558 2286 6634 2324
rect 6530 2226 6634 2286
rect 6530 2098 6604 2226
rect 6530 2078 6606 2098
rect 6586 2016 6676 2074
<< locali >>
rect 3714 2642 7904 2662
rect 3714 2576 3746 2642
rect 4110 2640 4384 2642
rect 4762 2640 5680 2642
rect 7872 2576 7904 2642
rect 3714 2468 7904 2576
rect 3714 2088 3942 2468
rect 7774 2088 7904 2468
rect 3714 2074 6612 2088
rect 6644 2074 7904 2088
rect 3714 1962 7904 2074
rect 3714 1960 7906 1962
rect 3714 1958 7904 1960
rect 41666 1474 41804 1478
rect 3348 856 41804 1474
rect 3348 408 3972 856
rect 5788 682 41804 856
rect 5788 664 8742 682
rect 8846 664 41804 682
rect 5788 662 6972 664
rect 7688 662 8742 664
rect 5788 408 6898 662
rect 3348 -158 6898 408
rect 7718 358 8742 662
rect 9590 458 10050 664
rect 10856 458 11316 664
rect 12162 458 12622 664
rect 13442 458 13902 664
rect 14734 458 15194 664
rect 16016 458 16476 664
rect 17326 656 41804 664
rect 17326 568 18496 656
rect 19332 568 19786 656
rect 20628 568 21050 656
rect 21920 568 22368 656
rect 23204 568 23650 656
rect 24472 568 24942 656
rect 25782 568 26236 656
rect 27022 654 41804 656
rect 17326 458 18504 568
rect 7710 -158 8742 358
rect 9574 -152 10054 458
rect 10856 284 11336 458
rect 10870 -152 11336 284
rect 12152 -152 12630 458
rect 13442 260 13920 458
rect 13446 -152 13920 260
rect 14732 -152 15200 458
rect 16008 -152 16482 458
rect 17308 -152 18504 458
rect 3348 -190 8742 -158
rect 8846 -158 18504 -152
rect 19318 512 19786 568
rect 19318 -158 19778 512
rect 20608 -158 21068 568
rect 21894 -158 22372 568
rect 23186 -158 23658 568
rect 24472 490 24948 568
rect 24482 -158 24948 490
rect 25760 512 26236 568
rect 25760 -158 26226 512
rect 27044 -158 41804 654
rect 8846 -190 41804 -158
rect 3348 -594 41804 -190
rect 3352 -608 41804 -594
rect 3352 -1364 3968 -608
rect 6436 -626 41804 -608
rect 34964 -1364 41804 -626
rect 3352 -1674 41804 -1364
rect 3348 -1728 41804 -1674
rect 3348 -9644 3974 -1728
rect 40466 -2368 41804 -1728
rect 40942 -9644 41804 -2368
rect 3348 -9804 41804 -9644
rect 3348 -9822 3430 -9804
rect 3350 -10040 3430 -9822
rect 41630 -10040 41804 -9804
rect 3350 -10156 41804 -10040
rect 40824 -10158 41804 -10156
rect 40824 -10160 41758 -10158
rect 40942 -10162 41758 -10160
<< viali >>
rect 3746 2640 4110 2642
rect 4384 2640 4762 2642
rect 5680 2640 7872 2642
rect 3746 2576 7872 2640
rect 3430 -10040 41630 -9804
<< metal1 >>
rect 3716 2642 7902 2662
rect 3716 2576 3746 2642
rect 4110 2640 4384 2642
rect 4762 2640 5680 2642
rect 7872 2576 7902 2642
rect 3716 2566 7902 2576
rect 3716 2554 7904 2566
rect 3718 2468 7904 2554
rect 3972 2460 4036 2468
rect 3972 2408 4032 2460
rect 3970 2396 4032 2408
rect 3970 2322 4030 2396
rect 4064 2358 4074 2410
rect 4408 2358 4418 2410
rect 4612 2398 4672 2468
rect 4610 2392 4672 2398
rect 3970 2234 4052 2322
rect 3986 2232 4052 2234
rect 4124 2154 4358 2358
rect 4436 2326 4470 2330
rect 4436 2260 4508 2326
rect 4610 2322 4670 2392
rect 4710 2362 4720 2414
rect 5054 2362 5064 2414
rect 5262 2400 5322 2468
rect 5260 2390 5322 2400
rect 4610 2308 4696 2322
rect 4436 2234 4510 2260
rect 4438 2232 4510 2234
rect 4454 2168 4510 2232
rect 4612 2232 4696 2308
rect 4612 2230 4672 2232
rect 4454 2040 4508 2168
rect 4770 2156 5004 2362
rect 5260 2324 5320 2390
rect 5360 2362 5370 2414
rect 5704 2362 5714 2414
rect 5260 2322 5324 2324
rect 5076 2314 5164 2320
rect 5076 2230 5114 2314
rect 5104 2138 5114 2230
rect 5172 2138 5182 2314
rect 5260 2234 5346 2322
rect 5286 2232 5346 2234
rect 5418 2154 5652 2362
rect 6008 2354 6018 2412
rect 6342 2354 6352 2412
rect 6654 2358 6664 2416
rect 6988 2358 6998 2416
rect 5906 2322 5974 2324
rect 5722 2320 5974 2322
rect 5722 2230 5988 2320
rect 5920 2226 5988 2230
rect 6072 2152 6290 2354
rect 6402 2320 6474 2324
rect 6558 2322 6634 2324
rect 6374 2238 6404 2320
rect 6394 2194 6404 2238
rect 6470 2194 6480 2320
rect 6534 2286 6634 2322
rect 6530 2226 6634 2286
rect 6402 2190 6474 2194
rect 5116 2096 5168 2138
rect 6530 2098 6604 2226
rect 6722 2152 6940 2358
rect 7290 2356 7300 2414
rect 7624 2356 7634 2414
rect 7018 2318 7090 2320
rect 7216 2318 7274 2322
rect 7018 2316 7106 2318
rect 7018 2238 7050 2316
rect 7034 2236 7050 2238
rect 7040 2174 7050 2236
rect 7114 2174 7124 2316
rect 7198 2226 7274 2318
rect 7198 2222 7262 2226
rect 7044 2170 7116 2174
rect 6530 2096 6612 2098
rect 5110 2040 6612 2096
rect 4452 2006 4534 2040
rect 6554 2038 6612 2040
rect 7200 2006 7262 2222
rect 7368 2154 7586 2356
rect 7660 2316 7732 2318
rect 7660 2236 7690 2316
rect 7680 2174 7690 2236
rect 7754 2174 7764 2316
rect 7684 2154 7756 2174
rect 4448 1956 7264 2006
rect 3560 1002 5370 1170
rect 3566 -708 3780 1002
rect 5302 870 5368 1002
rect 5302 862 5364 870
rect 5298 836 5364 862
rect 4026 708 4092 724
rect 4004 562 4014 708
rect 4082 562 4092 708
rect 4026 548 4092 562
rect 4146 512 4230 800
rect 4288 714 4336 718
rect 4288 711 4368 714
rect 4288 675 4447 711
rect 4287 543 4447 675
rect 4486 556 4496 728
rect 4550 556 4560 728
rect 4339 541 4447 543
rect 4502 546 4558 556
rect 4502 542 4556 546
rect 4066 450 4076 512
rect 4284 450 4294 512
rect 4397 295 4447 541
rect 4606 508 4690 796
rect 4748 552 5012 718
rect 4542 446 4552 508
rect 4760 446 4770 508
rect 5078 502 5162 798
rect 5298 712 5360 836
rect 5414 722 5460 724
rect 5216 706 5360 712
rect 5216 544 5366 706
rect 5398 536 5408 722
rect 5474 536 5484 722
rect 5000 450 5010 502
rect 5214 450 5224 502
rect 5410 295 5460 536
rect 5538 508 5622 792
rect 6084 714 6560 716
rect 5686 708 6560 714
rect 5686 540 6600 708
rect 8846 540 9020 582
rect 18606 558 19198 568
rect 19906 558 20498 568
rect 21196 558 21788 568
rect 22500 558 23092 568
rect 23758 558 24350 568
rect 25056 558 25648 568
rect 26350 560 26942 568
rect 26350 558 40155 560
rect 18580 552 40155 558
rect 18580 548 40892 552
rect 17164 540 17790 546
rect 5686 536 7604 540
rect 6084 528 7604 536
rect 5494 456 5504 508
rect 5708 456 5718 508
rect 4397 245 5460 295
rect 6290 -48 7604 528
rect 8846 526 17790 540
rect 8846 -38 17624 526
rect 8864 -44 17624 -38
rect 17164 -48 17624 -44
rect 6290 -50 6600 -48
rect 17614 -56 17624 -48
rect 17774 -48 17790 526
rect 17774 -56 17784 -48
rect 18580 -66 40944 548
rect 26364 -118 40944 -66
rect 27496 -170 40944 -118
rect 40058 -190 40944 -170
rect 3566 -1248 4466 -708
rect 35232 -758 35242 -752
rect 34472 -1280 35242 -758
rect 35232 -1300 35242 -1280
rect 35600 -758 35610 -752
rect 35600 -1280 35620 -758
rect 35600 -1300 35610 -1280
rect 4052 -3148 4460 -1836
rect 40466 -2368 40944 -190
rect 40466 -2384 40874 -2368
rect 4058 -4746 4466 -3434
rect 40456 -3968 40864 -2656
rect 4052 -6328 4460 -5016
rect 40472 -5550 40880 -4238
rect 4058 -7928 4466 -6616
rect 40458 -7138 40866 -5826
rect 4068 -9510 4476 -8198
rect 40464 -8754 40872 -7442
rect 40442 -8998 41668 -8974
rect 40442 -9536 41258 -8998
rect 41650 -9536 41668 -8998
rect 40442 -9540 41668 -9536
rect 3356 -9804 41748 -9648
rect 3356 -10040 3430 -9804
rect 41630 -10040 41748 -9804
rect 3356 -10162 41748 -10040
<< via1 >>
rect 4074 2358 4408 2410
rect 4720 2362 5054 2414
rect 5370 2362 5704 2414
rect 5114 2138 5172 2314
rect 6018 2354 6342 2412
rect 6664 2358 6988 2416
rect 6404 2194 6470 2320
rect 7300 2356 7624 2414
rect 7050 2174 7114 2316
rect 7690 2174 7754 2316
rect 4014 562 4082 708
rect 4496 556 4550 728
rect 4076 450 4284 512
rect 4552 446 4760 508
rect 5408 536 5474 722
rect 5010 450 5214 502
rect 5504 456 5708 508
rect 17624 -56 17774 526
rect 35242 -1300 35600 -752
rect 41258 -9536 41650 -8998
<< metal2 >>
rect 4762 2548 5018 2552
rect 5114 2548 5190 2552
rect 5410 2548 5666 2552
rect 4118 2476 5666 2548
rect 4118 2420 4374 2476
rect 4762 2424 5018 2476
rect 4074 2410 4408 2420
rect 4074 2348 4408 2358
rect 4720 2414 5054 2424
rect 4720 2352 5054 2362
rect 5114 2314 5190 2476
rect 5410 2424 5666 2476
rect 6064 2542 6318 2544
rect 6554 2542 6618 2544
rect 6688 2542 6942 2544
rect 7344 2542 7598 2544
rect 6064 2474 7598 2542
rect 5370 2414 5704 2424
rect 6064 2422 6318 2474
rect 6554 2460 6618 2474
rect 6688 2426 6942 2474
rect 5370 2352 5704 2362
rect 6018 2412 6342 2422
rect 6018 2344 6342 2354
rect 6664 2416 6988 2426
rect 6664 2348 6988 2358
rect 5172 2138 5190 2314
rect 6404 2327 6470 2330
rect 7082 2328 7180 2474
rect 7344 2424 7598 2474
rect 7300 2414 7624 2424
rect 7300 2346 7624 2356
rect 6404 2320 6522 2327
rect 7056 2326 7180 2328
rect 6470 2194 6522 2320
rect 6404 2184 6522 2194
rect 5114 2128 5190 2138
rect 6406 1907 6522 2184
rect 7050 2318 7180 2326
rect 7690 2322 7754 2326
rect 7050 2316 7188 2318
rect 7114 2174 7188 2316
rect 7050 2164 7188 2174
rect 3835 1759 6522 1907
rect 3835 1758 6470 1759
rect 3835 688 3936 1758
rect 7056 1648 7188 2164
rect 4390 1484 7188 1648
rect 7686 2316 7818 2322
rect 7686 2174 7690 2316
rect 7754 2174 7818 2316
rect 7686 1660 7818 2174
rect 40334 1660 40644 1664
rect 7686 1656 40862 1660
rect 41256 1656 41648 1658
rect 7686 1534 41648 1656
rect 7686 1528 40862 1534
rect 4390 728 4550 1484
rect 17780 1382 26068 1388
rect 17780 1374 28444 1382
rect 17780 974 35606 1374
rect 4014 708 4082 718
rect 3835 578 4014 688
rect 3835 277 3946 578
rect 4390 624 4496 728
rect 4392 592 4496 624
rect 4014 552 4082 562
rect 5408 722 5474 732
rect 4496 546 4550 556
rect 5382 536 5408 718
rect 17780 608 18186 974
rect 20156 968 35606 974
rect 27318 960 35606 968
rect 17736 536 18186 608
rect 5382 528 5474 536
rect 5386 526 5474 528
rect 17624 526 18186 536
rect 4076 512 4284 522
rect 4076 440 4284 450
rect 4552 508 4760 518
rect 4096 277 4268 440
rect 4552 436 4760 446
rect 5010 502 5214 512
rect 5010 440 5214 450
rect 4570 277 4742 436
rect 3835 254 4742 277
rect 3835 190 4744 254
rect 5040 228 5202 440
rect 5386 228 5462 526
rect 5504 508 5708 518
rect 5504 446 5708 456
rect 5530 228 5686 446
rect 3835 183 4735 190
rect 3872 182 3946 183
rect 5040 182 5686 228
rect 5042 170 5686 182
rect 17774 268 18186 526
rect 17774 -56 18162 268
rect 17624 -66 18162 -56
rect 17638 -70 18162 -66
rect 35236 -752 35600 960
rect 35236 -1300 35242 -752
rect 35242 -1310 35600 -1300
rect 41256 -8634 41648 1534
rect 41256 -8704 41652 -8634
rect 41260 -8998 41652 -8704
rect 41650 -9536 41652 -8998
rect 41260 -9538 41652 -9536
use sky130_fd_pr__pfet_01v8_lvt_2CMFLT  XM1
timestamp 1739201171
transform 1 0 4242 0 1 2278
box -376 -264 376 264
use sky130_fd_pr__nfet_01v8_lvt_S3357R  XM2
timestamp 1739201171
transform 1 0 5116 0 1 632
box -286 -300 286 300
use sky130_fd_pr__pfet_01v8_lvt_2CMFLT  XM3
timestamp 1739201171
transform 1 0 4888 0 1 2278
box -376 -264 376 264
use sky130_fd_pr__nfet_01v8_lvt_S3357R  XM4
timestamp 1739201171
transform 1 0 4184 0 1 632
box -286 -300 286 300
use sky130_fd_pr__pfet_01v8_lvt_2CMFLT  XM5
timestamp 1739201171
transform 1 0 6826 0 1 2278
box -376 -264 376 264
use sky130_fd_pr__pfet_01v8_lvt_2CMFLT  XM6
timestamp 1739201171
transform 1 0 7472 0 1 2278
box -376 -264 376 264
use sky130_fd_pr__pfet_01v8_lvt_2CMFLT  XM7
timestamp 1739201171
transform 1 0 6180 0 1 2278
box -376 -264 376 264
use sky130_fd_pr__pfet_01v8_lvt_2CMFLT  XM8
timestamp 1739201171
transform 1 0 5534 0 1 2278
box -376 -264 376 264
use sky130_fd_pr__nfet_01v8_lvt_S3357R  XM9
timestamp 1739201171
transform 1 0 5582 0 1 632
box -286 -300 286 300
use sky130_fd_pr__nfet_01v8_lvt_S3357R  XM10
timestamp 1739201171
transform 1 0 4650 0 1 632
box -286 -300 286 300
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ1 ~/pdk/sky130A/libs.ref/sky130_fd_pr/mag
array 0 6 1288 0 0 1288
timestamp 1704896540
transform 1 0 18240 0 1 -422
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2
array 0 6 1288 0 0 1288
timestamp 1704896540
transform 1 0 8500 0 1 -416
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ3
timestamp 1704896540
transform 1 0 6636 0 1 -418
box 0 0 1340 1340
use sky130_fd_pr__res_xhigh_po_2p85_FTTYMQ  XR2
timestamp 1739201171
transform 0 1 19470 -1 0 -987
box -451 -15582 451 15582
use sky130_fd_pr__res_xhigh_po_2p85_V69GM6  XR3
timestamp 1739201171
transform 0 1 22458 -1 0 -9271
box -451 -18582 451 18582
use sky130_fd_pr__res_xhigh_po_2p85_V69GM6  XR4
timestamp 1739201171
transform 0 1 22458 -1 0 -2107
box -451 -18582 451 18582
use sky130_fd_pr__res_xhigh_po_2p85_V69GM6  XR5
timestamp 1739201171
transform 0 1 22458 -1 0 -2903
box -451 -18582 451 18582
use sky130_fd_pr__res_xhigh_po_2p85_V69GM6  XR6
timestamp 1739201171
transform 0 1 22458 -1 0 -3699
box -451 -18582 451 18582
use sky130_fd_pr__res_xhigh_po_2p85_V69GM6  XR7
timestamp 1739201171
transform 0 -1 22458 1 0 -4495
box -451 -18582 451 18582
use sky130_fd_pr__res_xhigh_po_2p85_V69GM6  XR8
timestamp 1739201171
transform 0 1 22458 -1 0 -5291
box -451 -18582 451 18582
use sky130_fd_pr__res_xhigh_po_2p85_V69GM6  XR9
timestamp 1739201171
transform 0 1 22458 -1 0 -6087
box -451 -18582 451 18582
use sky130_fd_pr__res_xhigh_po_2p85_V69GM6  XR10
timestamp 1739201171
transform 0 1 22458 -1 0 -8475
box -451 -18582 451 18582
use sky130_fd_pr__res_xhigh_po_2p85_V69GM6  XR11
timestamp 1739201171
transform 0 1 22458 -1 0 -7679
box -451 -18582 451 18582
use sky130_fd_pr__res_xhigh_po_2p85_V69GM6  XR12
timestamp 1739201171
transform 0 1 22458 -1 0 -6883
box -451 -18582 451 18582
<< end >>
