MACRO bandgap
  CLASS BLOCK ;
  FOREIGN bandgap ;
  ORIGIN -16.740 50.810 ;
  SIZE 192.280 BY 64.120 ;
  OBS
      LAYER nwell ;
        RECT 19.330 10.070 39.240 12.710 ;
      LAYER pwell ;
        RECT 19.490 1.660 29.340 4.660 ;
        RECT 33.180 3.845 39.880 4.610 ;
        RECT 33.180 -1.325 33.945 3.845 ;
        RECT 39.115 -1.325 39.880 3.845 ;
        RECT 33.180 -2.090 39.880 -1.325 ;
        RECT 42.500 3.855 87.840 4.620 ;
        RECT 42.500 -1.315 43.265 3.855 ;
        RECT 48.435 -1.315 49.705 3.855 ;
        RECT 54.875 -1.315 56.145 3.855 ;
        RECT 61.315 -1.315 62.585 3.855 ;
        RECT 67.755 -1.315 69.025 3.855 ;
        RECT 74.195 -1.315 75.465 3.855 ;
        RECT 80.635 -1.315 81.905 3.855 ;
        RECT 87.075 -1.315 87.840 3.855 ;
        RECT 42.500 -2.080 87.840 -1.315 ;
        RECT 91.200 3.825 136.540 4.590 ;
        RECT 91.200 -1.345 91.965 3.825 ;
        RECT 97.135 -1.345 98.405 3.825 ;
        RECT 103.575 -1.345 104.845 3.825 ;
        RECT 110.015 -1.345 111.285 3.825 ;
        RECT 116.455 -1.345 117.725 3.825 ;
        RECT 122.895 -1.345 124.165 3.825 ;
        RECT 129.335 -1.345 130.605 3.825 ;
        RECT 135.775 -1.345 136.540 3.825 ;
        RECT 91.200 -2.110 136.540 -1.345 ;
        RECT 19.440 -7.190 175.260 -2.680 ;
        RECT 19.380 -48.610 205.200 -8.280 ;
      LAYER li1 ;
        RECT 18.570 12.340 39.520 13.310 ;
        RECT 18.570 10.440 19.710 12.340 ;
        RECT 20.310 11.850 22.110 12.020 ;
        RECT 20.080 11.145 20.250 11.635 ;
        RECT 22.170 11.145 22.340 11.635 ;
        RECT 20.310 10.760 22.110 10.930 ;
        RECT 22.740 10.440 22.910 12.340 ;
        RECT 23.540 11.850 25.340 12.020 ;
        RECT 23.310 11.145 23.480 11.635 ;
        RECT 25.400 11.145 25.570 11.635 ;
        RECT 23.540 10.760 25.340 10.930 ;
        RECT 25.970 10.440 26.140 12.340 ;
        RECT 26.770 11.850 28.570 12.020 ;
        RECT 26.540 11.145 26.710 11.635 ;
        RECT 28.630 11.145 28.800 11.635 ;
        RECT 26.770 10.760 28.570 10.930 ;
        RECT 29.200 10.440 29.370 12.340 ;
        RECT 30.000 11.850 31.800 12.020 ;
        RECT 29.770 11.145 29.940 11.635 ;
        RECT 31.860 11.145 32.030 11.635 ;
        RECT 30.000 10.760 31.800 10.930 ;
        RECT 32.430 10.440 32.600 12.340 ;
        RECT 33.230 11.850 35.030 12.020 ;
        RECT 33.000 11.145 33.170 11.635 ;
        RECT 35.090 11.145 35.260 11.635 ;
        RECT 33.230 10.760 35.030 10.930 ;
        RECT 35.660 10.440 35.830 12.340 ;
        RECT 36.460 11.850 38.260 12.020 ;
        RECT 36.230 11.145 36.400 11.635 ;
        RECT 38.320 11.145 38.490 11.635 ;
        RECT 36.460 10.760 38.260 10.930 ;
        RECT 38.870 10.440 39.520 12.340 ;
        RECT 18.570 9.790 39.520 10.440 ;
        RECT 208.330 7.370 209.020 7.390 ;
        RECT 16.740 4.280 209.020 7.370 ;
        RECT 16.740 2.040 19.860 4.280 ;
        RECT 20.470 3.800 21.370 3.970 ;
        RECT 20.240 2.690 20.410 3.630 ;
        RECT 21.430 2.690 21.600 3.630 ;
        RECT 20.470 2.350 21.370 2.520 ;
        RECT 22.000 2.040 22.170 4.280 ;
        RECT 22.800 3.800 23.700 3.970 ;
        RECT 22.570 2.690 22.740 3.630 ;
        RECT 23.760 2.690 23.930 3.630 ;
        RECT 22.800 2.350 23.700 2.520 ;
        RECT 24.330 2.040 24.500 4.280 ;
        RECT 25.130 3.800 26.030 3.970 ;
        RECT 24.900 2.690 25.070 3.630 ;
        RECT 26.090 2.690 26.260 3.630 ;
        RECT 25.130 2.350 26.030 2.520 ;
        RECT 26.660 2.040 26.830 4.280 ;
        RECT 27.460 3.800 28.360 3.970 ;
        RECT 27.230 2.690 27.400 3.630 ;
        RECT 28.420 2.690 28.590 3.630 ;
        RECT 28.940 3.315 209.020 4.280 ;
        RECT 28.940 3.305 43.805 3.315 ;
        RECT 27.460 2.350 28.360 2.520 ;
        RECT 28.940 2.040 34.490 3.305 ;
        RECT 16.740 -0.785 34.490 2.040 ;
        RECT 34.795 -0.475 38.265 2.995 ;
        RECT 38.575 1.790 43.805 3.305 ;
        RECT 38.550 -0.775 43.805 1.790 ;
        RECT 44.115 -0.465 47.585 3.005 ;
        RECT 47.895 2.290 50.250 3.315 ;
        RECT 47.870 -0.760 50.270 2.290 ;
        RECT 50.555 -0.465 54.025 3.005 ;
        RECT 54.280 1.420 56.685 3.315 ;
        RECT 54.335 -0.760 56.685 1.420 ;
        RECT 56.995 -0.465 60.465 3.005 ;
        RECT 60.775 2.290 63.125 3.315 ;
        RECT 60.760 -0.760 63.150 2.290 ;
        RECT 63.435 -0.465 66.905 3.005 ;
        RECT 67.210 2.290 69.565 3.315 ;
        RECT 67.210 1.300 69.600 2.290 ;
        RECT 67.215 -0.760 69.600 1.300 ;
        RECT 69.875 -0.465 73.345 3.005 ;
        RECT 73.655 -0.760 76.005 3.315 ;
        RECT 76.315 -0.465 79.785 3.005 ;
        RECT 80.080 2.290 82.445 3.315 ;
        RECT 86.535 3.280 209.020 3.315 ;
        RECT 80.040 -0.760 82.445 2.290 ;
        RECT 82.755 -0.465 86.225 3.005 ;
        RECT 86.535 2.840 92.505 3.280 ;
        RECT 86.535 -0.760 92.520 2.840 ;
        RECT 92.815 -0.495 96.285 2.975 ;
        RECT 96.595 2.840 98.945 3.280 ;
        RECT 44.230 -0.775 92.520 -0.760 ;
        RECT 38.550 -0.785 92.520 -0.775 ;
        RECT 16.740 -0.790 92.520 -0.785 ;
        RECT 96.590 -0.790 98.945 2.840 ;
        RECT 99.255 -0.495 102.725 2.975 ;
        RECT 103.035 -0.790 105.385 3.280 ;
        RECT 105.695 -0.495 109.165 2.975 ;
        RECT 109.475 2.840 111.840 3.280 ;
        RECT 109.470 -0.790 111.860 2.840 ;
        RECT 112.135 -0.495 115.605 2.975 ;
        RECT 115.915 2.840 118.265 3.280 ;
        RECT 115.915 -0.790 118.290 2.840 ;
        RECT 118.575 -0.495 122.045 2.975 ;
        RECT 122.355 2.840 124.710 3.280 ;
        RECT 122.355 -0.790 124.740 2.840 ;
        RECT 125.015 -0.495 128.485 2.975 ;
        RECT 128.795 2.560 131.180 3.280 ;
        RECT 135.110 3.270 209.020 3.280 ;
        RECT 128.795 -0.790 131.145 2.560 ;
        RECT 131.455 -0.495 134.925 2.975 ;
        RECT 135.220 -0.790 209.020 3.270 ;
        RECT 16.740 -2.970 209.020 -0.790 ;
        RECT 16.760 -3.040 209.020 -2.970 ;
        RECT 16.760 -6.820 19.840 -3.040 ;
        RECT 32.180 -3.130 209.020 -3.040 ;
        RECT 20.270 -6.360 22.430 -3.510 ;
        RECT 172.270 -6.360 174.430 -3.510 ;
        RECT 174.820 -6.820 209.020 -3.130 ;
        RECT 16.760 -8.370 209.020 -6.820 ;
        RECT 16.740 -8.640 209.020 -8.370 ;
        RECT 16.740 -12.440 19.870 -8.640 ;
        RECT 202.330 -9.110 209.020 -8.640 ;
        RECT 20.210 -11.960 22.370 -9.110 ;
        RECT 202.210 -11.840 209.020 -9.110 ;
        RECT 202.210 -11.960 204.370 -11.840 ;
        RECT 204.710 -12.440 209.020 -11.840 ;
        RECT 16.740 -12.610 209.020 -12.440 ;
        RECT 16.740 -16.420 19.870 -12.610 ;
        RECT 20.210 -15.940 22.370 -13.090 ;
        RECT 202.210 -15.940 204.370 -13.090 ;
        RECT 204.710 -16.420 209.020 -12.610 ;
        RECT 16.740 -16.590 209.020 -16.420 ;
        RECT 16.740 -20.400 19.870 -16.590 ;
        RECT 20.210 -19.920 22.370 -17.070 ;
        RECT 202.210 -19.920 204.370 -17.070 ;
        RECT 204.710 -20.400 209.020 -16.590 ;
        RECT 16.740 -20.570 209.020 -20.400 ;
        RECT 16.740 -24.380 19.870 -20.570 ;
        RECT 20.210 -23.900 22.370 -21.050 ;
        RECT 202.210 -23.900 204.370 -21.050 ;
        RECT 204.710 -24.380 209.020 -20.570 ;
        RECT 16.740 -24.550 209.020 -24.380 ;
        RECT 16.740 -28.360 19.870 -24.550 ;
        RECT 20.210 -27.880 22.370 -25.030 ;
        RECT 202.210 -27.880 204.370 -25.030 ;
        RECT 204.710 -28.360 209.020 -24.550 ;
        RECT 16.740 -28.530 209.020 -28.360 ;
        RECT 16.740 -32.340 19.870 -28.530 ;
        RECT 20.210 -31.860 22.370 -29.010 ;
        RECT 202.210 -31.860 204.370 -29.010 ;
        RECT 204.710 -32.340 209.020 -28.530 ;
        RECT 16.740 -32.510 209.020 -32.340 ;
        RECT 16.740 -36.320 19.870 -32.510 ;
        RECT 20.210 -35.840 22.370 -32.990 ;
        RECT 202.210 -35.840 204.370 -32.990 ;
        RECT 204.710 -36.320 209.020 -32.510 ;
        RECT 16.740 -36.490 209.020 -36.320 ;
        RECT 16.740 -40.300 19.870 -36.490 ;
        RECT 20.210 -39.820 22.370 -36.970 ;
        RECT 202.210 -39.820 204.370 -36.970 ;
        RECT 204.710 -40.300 209.020 -36.490 ;
        RECT 16.740 -40.470 209.020 -40.300 ;
        RECT 16.740 -44.280 19.870 -40.470 ;
        RECT 20.210 -43.800 22.370 -40.950 ;
        RECT 202.210 -43.800 204.370 -40.950 ;
        RECT 204.710 -44.280 209.020 -40.470 ;
        RECT 16.740 -44.450 209.020 -44.280 ;
        RECT 16.740 -48.220 19.870 -44.450 ;
        RECT 20.210 -47.780 22.370 -44.930 ;
        RECT 202.210 -47.780 204.370 -44.930 ;
        RECT 204.710 -48.220 209.020 -44.450 ;
        RECT 16.740 -49.110 209.020 -48.220 ;
        RECT 16.750 -50.780 209.020 -49.110 ;
        RECT 204.120 -50.790 209.020 -50.780 ;
        RECT 204.120 -50.800 208.790 -50.790 ;
        RECT 204.710 -50.810 208.790 -50.800 ;
      LAYER met1 ;
        RECT 18.580 12.830 39.510 13.310 ;
        RECT 18.580 12.770 39.520 12.830 ;
        RECT 18.590 12.340 39.520 12.770 ;
        RECT 19.860 12.300 20.180 12.340 ;
        RECT 19.860 12.040 20.160 12.300 ;
        RECT 19.850 11.980 20.160 12.040 ;
        RECT 19.850 11.615 20.150 11.980 ;
        RECT 20.320 11.790 22.090 12.050 ;
        RECT 23.060 11.990 23.360 12.340 ;
        RECT 23.050 11.960 23.360 11.990 ;
        RECT 19.850 11.170 20.280 11.615 ;
        RECT 19.930 11.165 20.280 11.170 ;
        RECT 19.930 11.160 20.260 11.165 ;
        RECT 20.620 10.960 21.790 11.790 ;
        RECT 22.180 11.630 22.350 11.650 ;
        RECT 22.180 11.615 22.540 11.630 ;
        RECT 22.140 11.300 22.540 11.615 ;
        RECT 23.050 11.615 23.350 11.960 ;
        RECT 23.550 11.810 25.320 12.070 ;
        RECT 26.310 12.000 26.610 12.340 ;
        RECT 26.800 12.050 28.570 12.070 ;
        RECT 30.040 12.050 31.760 12.060 ;
        RECT 33.270 12.050 34.990 12.080 ;
        RECT 36.450 12.050 38.170 12.070 ;
        RECT 26.300 11.950 26.610 12.000 ;
        RECT 23.050 11.540 23.510 11.615 ;
        RECT 22.140 11.165 22.550 11.300 ;
        RECT 22.190 11.160 22.550 11.165 ;
        RECT 20.330 10.730 22.090 10.960 ;
        RECT 22.270 10.840 22.550 11.160 ;
        RECT 23.060 11.165 23.510 11.540 ;
        RECT 23.060 11.160 23.480 11.165 ;
        RECT 23.060 11.150 23.360 11.160 ;
        RECT 23.850 10.960 25.020 11.810 ;
        RECT 26.300 11.620 26.600 11.950 ;
        RECT 26.790 11.820 28.570 12.050 ;
        RECT 30.020 11.820 31.780 12.050 ;
        RECT 33.250 11.820 35.010 12.050 ;
        RECT 36.450 11.820 38.240 12.050 ;
        RECT 26.800 11.810 28.570 11.820 ;
        RECT 26.300 11.615 26.620 11.620 ;
        RECT 25.370 11.600 25.600 11.615 ;
        RECT 25.370 11.570 25.820 11.600 ;
        RECT 25.370 11.165 25.910 11.570 ;
        RECT 26.300 11.170 26.740 11.615 ;
        RECT 25.380 11.150 25.910 11.165 ;
        RECT 26.430 11.165 26.740 11.170 ;
        RECT 26.430 11.160 26.730 11.165 ;
        RECT 22.270 10.200 22.540 10.840 ;
        RECT 23.560 10.730 25.320 10.960 ;
        RECT 25.520 10.690 25.910 11.150 ;
        RECT 27.090 10.960 28.260 11.810 ;
        RECT 30.040 11.770 31.760 11.820 ;
        RECT 33.270 11.790 34.990 11.820 ;
        RECT 29.530 11.615 29.870 11.620 ;
        RECT 28.600 11.610 28.830 11.615 ;
        RECT 29.530 11.610 29.970 11.615 ;
        RECT 28.600 11.165 29.970 11.610 ;
        RECT 28.610 11.150 29.940 11.165 ;
        RECT 29.600 11.130 29.940 11.150 ;
        RECT 30.360 10.960 31.450 11.770 ;
        RECT 32.010 11.615 32.370 11.620 ;
        RECT 31.830 11.600 32.370 11.615 ;
        RECT 32.790 11.615 33.170 11.620 ;
        RECT 32.790 11.610 33.200 11.615 ;
        RECT 31.830 11.165 32.400 11.600 ;
        RECT 32.670 11.430 33.200 11.610 ;
        RECT 31.970 10.970 32.400 11.165 ;
        RECT 32.650 11.165 33.200 11.430 ;
        RECT 32.650 11.130 33.170 11.165 ;
        RECT 26.790 10.730 28.550 10.960 ;
        RECT 30.020 10.730 31.780 10.960 ;
        RECT 32.010 10.950 32.370 10.970 ;
        RECT 25.580 10.480 25.840 10.690 ;
        RECT 32.650 10.490 33.020 11.130 ;
        RECT 33.610 10.960 34.700 11.790 ;
        RECT 36.450 11.780 38.170 11.820 ;
        RECT 35.060 11.600 35.290 11.615 ;
        RECT 36.200 11.610 36.430 11.615 ;
        RECT 35.060 11.590 35.450 11.600 ;
        RECT 36.080 11.590 36.430 11.610 ;
        RECT 35.060 11.580 35.530 11.590 ;
        RECT 35.060 11.165 35.620 11.580 ;
        RECT 33.250 10.730 35.010 10.960 ;
        RECT 35.200 10.870 35.620 11.165 ;
        RECT 35.990 11.165 36.430 11.590 ;
        RECT 35.990 11.130 36.370 11.165 ;
        RECT 35.990 11.110 36.310 11.130 ;
        RECT 35.220 10.850 35.580 10.870 ;
        RECT 32.650 10.480 33.060 10.490 ;
        RECT 25.550 10.200 33.060 10.480 ;
        RECT 22.260 10.030 22.670 10.200 ;
        RECT 32.770 10.190 33.060 10.200 ;
        RECT 36.000 10.030 36.310 11.110 ;
        RECT 36.840 10.960 37.930 11.780 ;
        RECT 38.290 11.590 38.520 11.615 ;
        RECT 38.290 11.580 38.660 11.590 ;
        RECT 38.290 11.165 38.820 11.580 ;
        RECT 36.480 10.730 38.240 10.960 ;
        RECT 38.400 10.870 38.820 11.165 ;
        RECT 38.420 10.770 38.780 10.870 ;
        RECT 22.240 9.780 36.320 10.030 ;
        RECT 17.800 5.010 26.850 5.850 ;
        RECT 17.830 -3.540 18.900 5.010 ;
        RECT 26.510 4.350 26.840 5.010 ;
        RECT 26.510 4.310 26.820 4.350 ;
        RECT 26.490 4.180 26.820 4.310 ;
        RECT 20.490 3.770 21.350 4.000 ;
        RECT 22.820 3.770 23.680 4.000 ;
        RECT 25.150 3.770 26.010 4.000 ;
        RECT 20.130 3.540 20.460 3.620 ;
        RECT 20.020 2.810 20.460 3.540 ;
        RECT 20.130 2.740 20.460 2.810 ;
        RECT 20.210 2.710 20.440 2.740 ;
        RECT 20.730 2.560 21.150 3.770 ;
        RECT 21.400 3.590 21.630 3.610 ;
        RECT 21.400 3.570 21.680 3.590 ;
        RECT 21.400 3.555 21.840 3.570 ;
        RECT 21.400 2.710 22.180 3.555 ;
        RECT 22.540 3.530 22.770 3.610 ;
        RECT 22.360 2.980 22.790 3.530 ;
        RECT 22.540 2.710 22.770 2.980 ;
        RECT 21.550 2.705 22.180 2.710 ;
        RECT 21.550 2.700 21.810 2.705 ;
        RECT 20.330 2.250 21.470 2.560 ;
        RECT 21.985 2.050 22.180 2.705 ;
        RECT 23.050 2.550 23.430 3.770 ;
        RECT 23.730 3.590 23.960 3.610 ;
        RECT 24.870 3.590 25.100 3.610 ;
        RECT 23.730 2.770 25.100 3.590 ;
        RECT 23.730 2.710 23.960 2.770 ;
        RECT 24.140 2.760 25.100 2.770 ;
        RECT 24.870 2.710 25.100 2.760 ;
        RECT 25.390 2.550 25.810 3.770 ;
        RECT 26.060 3.560 26.290 3.610 ;
        RECT 26.490 3.560 26.800 4.180 ;
        RECT 27.480 3.770 28.340 4.000 ;
        RECT 27.070 3.610 27.300 3.620 ;
        RECT 26.060 3.530 26.800 3.560 ;
        RECT 26.060 2.720 26.830 3.530 ;
        RECT 26.060 2.710 26.290 2.720 ;
        RECT 26.990 2.710 27.430 3.610 ;
        RECT 26.990 2.680 27.420 2.710 ;
        RECT 22.820 2.510 23.680 2.550 ;
        RECT 25.150 2.510 26.010 2.550 ;
        RECT 22.810 2.220 23.690 2.510 ;
        RECT 25.000 2.250 26.120 2.510 ;
        RECT 21.985 1.475 22.235 2.050 ;
        RECT 27.050 1.475 27.300 2.680 ;
        RECT 27.690 2.550 28.110 3.770 ;
        RECT 28.390 3.570 28.620 3.610 ;
        RECT 30.420 3.570 32.800 3.580 ;
        RECT 28.390 3.540 32.800 3.570 ;
        RECT 28.390 2.710 33.000 3.540 ;
        RECT 44.230 2.795 45.100 2.910 ;
        RECT 28.430 2.700 33.000 2.710 ;
        RECT 35.005 2.700 38.055 2.785 ;
        RECT 28.430 2.680 38.055 2.700 ;
        RECT 30.420 2.640 38.055 2.680 ;
        RECT 27.480 2.540 28.340 2.550 ;
        RECT 27.470 2.280 28.590 2.540 ;
        RECT 21.985 1.225 27.300 1.475 ;
        RECT 31.450 -0.240 38.055 2.640 ;
        RECT 44.230 2.700 47.375 2.795 ;
        RECT 50.765 2.700 53.815 2.795 ;
        RECT 57.205 2.700 60.255 2.795 ;
        RECT 63.645 2.700 66.695 2.795 ;
        RECT 70.085 2.700 73.135 2.795 ;
        RECT 76.525 2.700 79.575 2.795 ;
        RECT 82.965 2.730 86.015 2.795 ;
        RECT 93.030 2.790 95.990 2.840 ;
        RECT 99.530 2.790 102.490 2.840 ;
        RECT 105.980 2.790 108.940 2.840 ;
        RECT 112.500 2.790 115.460 2.840 ;
        RECT 118.790 2.790 121.750 2.840 ;
        RECT 125.280 2.790 128.240 2.840 ;
        RECT 131.750 2.800 134.710 2.840 ;
        RECT 131.750 2.790 200.775 2.800 ;
        RECT 92.900 2.760 200.775 2.790 ;
        RECT 92.900 2.740 204.460 2.760 ;
        RECT 82.965 2.700 88.950 2.730 ;
        RECT 44.230 -0.190 88.950 2.700 ;
        RECT 44.320 -0.220 88.950 -0.190 ;
        RECT 31.450 -0.250 33.000 -0.240 ;
        RECT 35.005 -0.265 38.055 -0.240 ;
        RECT 44.325 -0.255 47.375 -0.220 ;
        RECT 50.765 -0.255 53.815 -0.220 ;
        RECT 57.205 -0.255 60.255 -0.220 ;
        RECT 63.645 -0.255 66.695 -0.220 ;
        RECT 70.085 -0.255 73.135 -0.220 ;
        RECT 76.525 -0.255 79.575 -0.220 ;
        RECT 82.965 -0.240 88.950 -0.220 ;
        RECT 82.965 -0.255 86.015 -0.240 ;
        RECT 88.070 -0.280 88.920 -0.240 ;
        RECT 92.900 -0.330 204.720 2.740 ;
        RECT 131.820 -0.590 204.720 -0.330 ;
        RECT 137.480 -0.850 204.720 -0.590 ;
        RECT 200.290 -0.950 204.720 -0.850 ;
        RECT 20.330 -3.540 22.375 -3.530 ;
        RECT 17.830 -6.240 22.375 -3.540 ;
        RECT 20.330 -6.340 22.375 -6.240 ;
        RECT 172.325 -3.790 174.370 -3.530 ;
        RECT 176.160 -3.790 178.050 -3.760 ;
        RECT 172.325 -6.340 178.100 -3.790 ;
        RECT 172.360 -6.400 178.100 -6.340 ;
        RECT 176.160 -6.500 178.050 -6.400 ;
        RECT 202.330 -9.130 204.720 -0.950 ;
        RECT 20.270 -9.180 22.315 -9.130 ;
        RECT 20.260 -11.940 22.315 -9.180 ;
        RECT 202.265 -11.840 204.720 -9.130 ;
        RECT 202.265 -11.920 204.370 -11.840 ;
        RECT 202.265 -11.940 204.310 -11.920 ;
        RECT 20.260 -13.110 22.300 -11.940 ;
        RECT 20.260 -15.740 22.315 -13.110 ;
        RECT 20.270 -15.920 22.315 -15.740 ;
        RECT 202.265 -13.280 204.310 -13.110 ;
        RECT 202.265 -15.920 204.320 -13.280 ;
        RECT 202.280 -17.090 204.320 -15.920 ;
        RECT 20.270 -17.170 22.315 -17.090 ;
        RECT 20.270 -19.900 22.330 -17.170 ;
        RECT 202.265 -19.840 204.320 -17.090 ;
        RECT 202.265 -19.900 204.310 -19.840 ;
        RECT 20.290 -21.070 22.330 -19.900 ;
        RECT 20.270 -23.730 22.330 -21.070 ;
        RECT 202.265 -21.190 204.310 -21.070 ;
        RECT 20.270 -23.880 22.315 -23.730 ;
        RECT 202.265 -23.880 204.400 -21.190 ;
        RECT 202.360 -25.050 204.400 -23.880 ;
        RECT 20.270 -25.080 22.315 -25.050 ;
        RECT 20.260 -27.860 22.315 -25.080 ;
        RECT 202.265 -27.750 204.400 -25.050 ;
        RECT 202.265 -27.860 204.310 -27.750 ;
        RECT 20.260 -29.030 22.300 -27.860 ;
        RECT 20.260 -31.640 22.315 -29.030 ;
        RECT 20.270 -31.840 22.315 -31.640 ;
        RECT 202.265 -29.130 204.310 -29.030 ;
        RECT 202.265 -31.840 204.330 -29.130 ;
        RECT 202.290 -33.010 204.330 -31.840 ;
        RECT 20.270 -33.080 22.315 -33.010 ;
        RECT 20.270 -35.820 22.330 -33.080 ;
        RECT 202.265 -35.690 204.330 -33.010 ;
        RECT 202.265 -35.820 204.310 -35.690 ;
        RECT 20.290 -36.990 22.330 -35.820 ;
        RECT 20.270 -39.640 22.330 -36.990 ;
        RECT 202.265 -37.210 204.310 -36.990 ;
        RECT 20.270 -39.800 22.315 -39.640 ;
        RECT 202.265 -39.800 204.360 -37.210 ;
        RECT 202.320 -40.970 204.360 -39.800 ;
        RECT 20.270 -40.990 22.315 -40.970 ;
        RECT 20.270 -43.780 22.380 -40.990 ;
        RECT 202.265 -43.770 204.360 -40.970 ;
        RECT 202.265 -43.780 204.310 -43.770 ;
        RECT 20.340 -44.950 22.380 -43.780 ;
        RECT 206.100 -44.870 208.140 -44.860 ;
        RECT 20.270 -47.550 22.380 -44.950 ;
        RECT 20.270 -47.760 22.315 -47.550 ;
        RECT 202.210 -47.700 208.140 -44.870 ;
        RECT 202.265 -47.760 204.310 -47.700 ;
        RECT 16.780 -50.810 208.740 -48.240 ;
      LAYER met2 ;
        RECT 23.810 12.740 25.090 12.760 ;
        RECT 25.570 12.740 25.950 12.760 ;
        RECT 27.050 12.740 28.330 12.760 ;
        RECT 20.590 12.380 28.330 12.740 ;
        RECT 20.590 12.100 21.870 12.380 ;
        RECT 23.810 12.120 25.090 12.380 ;
        RECT 20.370 11.740 22.040 12.100 ;
        RECT 23.600 11.760 25.270 12.120 ;
        RECT 25.570 10.640 25.950 12.380 ;
        RECT 27.050 12.120 28.330 12.380 ;
        RECT 30.320 12.710 31.590 12.720 ;
        RECT 32.770 12.710 33.090 12.720 ;
        RECT 33.440 12.710 34.710 12.720 ;
        RECT 36.720 12.710 37.990 12.720 ;
        RECT 30.320 12.370 37.990 12.710 ;
        RECT 26.850 11.760 28.520 12.120 ;
        RECT 30.320 12.110 31.590 12.370 ;
        RECT 33.440 12.130 34.710 12.370 ;
        RECT 30.090 11.720 31.710 12.110 ;
        RECT 33.320 11.740 34.940 12.130 ;
        RECT 32.020 11.635 32.350 11.650 ;
        RECT 35.410 11.640 35.900 12.370 ;
        RECT 36.720 12.120 37.990 12.370 ;
        RECT 36.500 11.730 38.120 12.120 ;
        RECT 32.020 10.920 32.610 11.635 ;
        RECT 35.280 11.630 35.900 11.640 ;
        RECT 32.030 9.535 32.610 10.920 ;
        RECT 35.250 11.590 35.900 11.630 ;
        RECT 38.450 11.610 38.770 11.630 ;
        RECT 35.250 10.820 35.940 11.590 ;
        RECT 19.175 8.795 32.610 9.535 ;
        RECT 19.175 8.790 32.350 8.795 ;
        RECT 19.175 3.440 19.680 8.790 ;
        RECT 35.280 8.240 35.940 10.820 ;
        RECT 21.950 7.420 35.940 8.240 ;
        RECT 38.430 8.300 39.090 11.610 ;
        RECT 201.670 8.300 203.220 8.320 ;
        RECT 38.430 8.280 204.310 8.300 ;
        RECT 206.280 8.280 208.240 8.290 ;
        RECT 38.430 7.670 208.240 8.280 ;
        RECT 38.430 7.640 204.310 7.670 ;
        RECT 21.950 4.270 22.750 7.420 ;
        RECT 88.900 6.910 130.340 6.940 ;
        RECT 88.900 6.870 142.220 6.910 ;
        RECT 88.900 4.870 178.030 6.870 ;
        RECT 21.950 3.610 22.540 4.270 ;
        RECT 20.070 3.440 20.410 3.590 ;
        RECT 19.175 2.890 20.410 3.440 ;
        RECT 21.950 3.580 22.550 3.610 ;
        RECT 27.040 3.590 27.370 3.660 ;
        RECT 21.950 3.120 22.740 3.580 ;
        RECT 21.960 2.960 22.740 3.120 ;
        RECT 22.130 2.950 22.740 2.960 ;
        RECT 22.410 2.930 22.740 2.950 ;
        RECT 19.175 1.385 19.730 2.890 ;
        RECT 20.070 2.760 20.410 2.890 ;
        RECT 26.910 2.640 27.370 3.590 ;
        RECT 88.900 3.040 90.930 4.870 ;
        RECT 100.780 4.840 178.030 4.870 ;
        RECT 136.590 4.800 178.030 4.840 ;
        RECT 88.680 2.680 90.930 3.040 ;
        RECT 26.930 2.630 27.370 2.640 ;
        RECT 20.380 2.200 21.420 2.610 ;
        RECT 22.860 2.290 23.640 2.560 ;
        RECT 20.480 1.385 21.340 2.200 ;
        RECT 22.850 1.385 23.710 2.290 ;
        RECT 25.050 2.200 26.070 2.560 ;
        RECT 19.175 1.270 23.710 1.385 ;
        RECT 19.175 0.950 23.720 1.270 ;
        RECT 25.200 1.140 26.010 2.200 ;
        RECT 26.930 1.140 27.310 2.630 ;
        RECT 27.520 2.230 28.540 2.590 ;
        RECT 27.650 1.140 28.430 2.230 ;
        RECT 19.175 0.915 23.675 0.950 ;
        RECT 19.360 0.910 19.730 0.915 ;
        RECT 25.200 0.910 28.430 1.140 ;
        RECT 25.210 0.850 28.430 0.910 ;
        RECT 88.120 1.340 90.930 2.680 ;
        RECT 88.120 -0.330 90.810 1.340 ;
        RECT 88.190 -0.350 90.810 -0.330 ;
        RECT 176.180 -6.500 178.000 4.800 ;
        RECT 176.210 -6.550 178.000 -6.500 ;
        RECT 206.280 -43.170 208.240 7.670 ;
        RECT 206.280 -43.520 208.260 -43.170 ;
        RECT 206.300 -44.630 208.260 -43.520 ;
        RECT 206.290 -44.730 208.260 -44.630 ;
        RECT 206.290 -46.410 208.240 -44.730 ;
        RECT 206.300 -47.710 208.240 -46.410 ;
  END
END bandgap
END LIBRARY

